module Test_FSM;




endmodule
